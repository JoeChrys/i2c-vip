
//`include "uvm_pkg.sv"
`include "uvm_macros.svh" 
`include "i2c_pkg.sv"
package i2c_test_pkg;

import uvm_pkg::*;
import i2c_pkg::*;

// * * * You can include different sequences for specific test bellow * * *

endpackage 

//------------------------------------------------------------------------------------------------------------


